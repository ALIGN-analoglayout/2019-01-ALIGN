VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO Switch_PMOS_10_1x1
  ORIGIN 0 0 ;
  FOREIGN Switch_PMOS_10_1x1 0 0 ;
  SIZE 0.432 BY 0.378 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.064 0.432 0.082 ;
    END
  END S
 
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.128 0.432 0.146 ;
    END
  END D
  
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
    END
  END D
END Switch_PMOS_10_1x1

MACRO Switch_NMOS_10_1x1
  ORIGIN 0 0 ;
  FOREIGN Switch_NMOS_10_1x1 0 0 ;
  SIZE 0.432 BY 0.378 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.064 0.432 0.082 ;
    END
  END S
 
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.128 0.432 0.146 ;
    END
  END D
  
  PIN G
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0 0.432 0.018 ;
    END
  END D
END Switch_NMOS_10_1x1

