MACRO SCM_NMOS
MACRO CMC_PMOS
MACRO CMC_NMOS
MACRO DP_NMOS
END LIBRARY
