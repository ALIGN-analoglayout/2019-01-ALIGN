VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO res_3.8K
  ORIGIN 0 0 ;
  FOREIGN res_3.8K 0 0 ;
  SIZE 2.034 BY 1 ;
  PIN LEFT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.018 0.018 ;
    END
  END LEFT
  PIN RIGHT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 2.016 0 2.034 0.018 ;
    END
  END RIGHT
  OBS
      LAYER M1 ;
        RECT 0.018 0.018 2.016 1 ;
      END
END res_3.8K

MACRO res_3K
  ORIGIN 0 0 ;
  FOREIGN res_3K 0 0 ;
  SIZE 1.602 BY 1 ;
  PIN LEFT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0 0 0.018 0.018 ;
    END
  END LEFT
  PIN RIGHT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.584 0 1.602 0.018 ;
    END
  END RIGHT
  OBS
      LAYER M1 ;
        RECT 0.018 0.018 1.584 1 ;
      END
END res_3K

MACRO DP_NMOS_2x2_4x3
  ORIGIN 0 0 ;
  FOREIGN DP_NMOS_2x2_4x3 0 0 ;
  SIZE 0.864 BY 0.864 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.064 0.864 0.082 ;
    END
  END S
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.192 0.864 0.210 ;
    END
  END D1
  
  PIN D2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.128 0.864 0.146 ;
    END
  END D2

PIN G1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0 0.864 0.018 ;
    END
  END G1

PIN G2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.256 0.864 0.274 ;
    END
  END G2
 
  
END DP_NMOS_2x2_4x3

MACRO SCM_NMOS_4x4_4x3
  ORIGIN 0 0 ;
  FOREIGN SCM_NMOS_4x4_4x3 0 0 ;
  SIZE 0.864 BY 1.728 ;
  PIN S
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.064 0.864 0.082 ;
    END
  END S
  PIN D1
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.192 0.864 0.210 ;
    END
  END D1
  
  PIN D2
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0 0.128 0.864 0.146 ;
    END
  END D2
 
  
END SCM_NMOS_4x4_4x3

